-------------------------------------------------------
-- uProgramMemory
-- Cristian Durán
--	Organización de computadores
--	06-06-2022
-------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
-----------------------------------------------------
ENTITY uProgramMemory IS
PORT(	
		uaddr	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
		U_I	: 	OUT 	STD_LOGIC_VECTOR(28 DOWNTO 0));
END ENTITY uProgramMemory;
-----------------------------------------------------
ARCHITECTURE behavioral OF uProgramMemory IS
BEGIN
	
	MU_I: PROCESS(uaddr) 
	BEGIN
		CASE uaddr IS
	-- Complete the following values according to your particular implementation 
	-- Unused postions do not affect the operation of the ROM
			-- FETCH 							    
			WHEN "00000000" => U_I <= "00000000000100000000010110100"; 
			WHEN "00000001" => U_I <= "00000010000000000000010000000"; 
			WHEN "00000010" => U_I <= "00110001000000010000010000000"; 
			WHEN "00000011" => U_I <= "00000100000000100000001000000"; 
																					
			-- INT
			WHEN "00000100" => U_I <= "00000000000000000000110000000"; 
			WHEN "00000101" => U_I <= "00000000000000000000000000000"; 
			WHEN "00000110" => U_I <= "00000000000000000000000000000"; 
			WHEN "00000111" => U_I <= "00000000000000000000000000000"; 

			--00001	 MOV ACC,A 
			WHEN "00001000" => U_I <= "00000001111011000101001000000";
         WHEN "00001001" => U_I <= "00000000000000000000000000000";
			WHEN "00001010" => U_I <= "00000000000000000000000000000";
			WHEN "00001011" => U_I <= "00000000000000000000000000000";
			WHEN "00001100" => U_I <= "00000000000000000000000000000";
			WHEN "00001101" => U_I <= "00000000000000000000000000000";
			WHEN "00001110" => U_I <= "00000000000000000000000000000";  
			WHEN "00001111" => U_I <= "00000000000000000000000000000";
			
			
			
			--00010  MOV A,ACC
			WHEN "00010000" => U_I <= "00000001011111000101111000000";
			when "00010001" => U_I <= "00000000000000000000000000000";
			when "00010010" => U_I <= "00000000000000000000000000000";
			when "00010011" => U_I <= "00000000000000000000000000000";
			when "00010100" => U_I <= "00000000000000000000000000000";
			when "00010101" => U_I <= "00000000000000000000000000000";
			when "00010110" => U_I <= "00000000000000000000000000000";
			when "00010111" => U_I <= "00000000000000000000000000000";
			
			
			--00011	 MOV ACC,CTE
			WHEN "00011000" => U_I <= "00000010000000000000010000000";
			WHEN "00011001" => U_I <= "00110001000000010000010000000";
			WHEN "00011010" => U_I <= "00000001111000100001001000000";
         WHEN "00011011" => U_I <=  "00000000000000000000000000000";
			
			--00100  MOV ACC,[DPTR]
			WHEN "00100000" => U_I <= "00000010000010000000010000000";
			WHEN "00100001" => U_I <= "00000000000000110000010000000";
			WHEN "00100010" => U_I <= "00000001111000100001001000000";

			--00101  MOV DPTR,ACC
			WHEN "00101000" => U_I <= "00000001010111000100000000000";
			WHEN "00101001" => U_I <=  "00000000000000000000000000000";
			
			-- 00110 MOV [DPTR],ACC	
			WHEN "00110000" => U_I <= "00000010000010000011101000000";
			WHEN "00110001" => U_I <= "00000001001111101110000000000";
			WHEN "00110010" => U_I  <= "00000000000000000000000000000";	  
			

			-- 00111 INV ACC
			WHEN "00111000" => U_I <= "00001010000000000100000000000";
			WHEN "00111001" => U_I <=  "00000000000000000000000000000";	
			 -- 01000 AND ACC,A	 
			WHEN "01000000" => U_I <= "00000001010100000100000000000";
         WHEN "01000001" => U_I <=  "00000000000000000000000000000"; -- 
			
			-- 01001 ADD ACC,A
			WHEN "01001000" => U_I <= "00101001111011000100000000000";
			when "01001001" => U_I <=  "00000000000000000000000000000";
			
			-- 01010 JMP DIR
			WHEN "01010000" => U_I <= "00000010000000000011111001000";
			WHEN "01010001" => U_I <= "00110001000000010011111000000";
			WHEN "01010010" => U_I <= "00000010001000000010000000000";
			WHEN "01010011" => U_I <=  "00000000000000000000000000000";
			
			-- 01011 JZ DIR
			WHEN "01011000" => U_I <= "00000000000000000001111001000";
			WHEN "01011001" => U_I <= "00000001010000000000000000000";
			WHEN "01011010" => U_I <= "00000010000010000011111000000";
			WHEN "01011011" => U_I <= "00000100001000110010000000000";
			WHEN "01011100" => U_I <= "00000000000000000000000000000"; 
			
			-- 01100 JN DIR
			WHEN "01100000" => U_I <= "00000000000000000001111011000";
			WHEN "01100001" => U_I <= "00000100000000100000001000000";
			WHEN "01100010" => U_I <= "00000010000001000011111000000";
			WHEN "01100011" => U_I <= "00000100001000110010000000000";
			WHEN "01100100" => U_I <=  "00000000000000000000000000000";
			
			-- 01101 JC DIR
			WHEN "01101000" => U_I <= "00000000000000000000010100010";
			WHEN "01101001" => U_I <= "00110001000000000001000000000";
			WHEN "01101010" => U_I <= "00000010000000000000010000000";
			WHEN "01101011" => U_I <= "00000000000000110000010000000";
			WHEN "01101100" => U_I <= "00000001000000010001001000000";
			
			
			-- 01110  CALL DIR       
			WHEN "01110000" => U_I <= "00000010000001000011111000000";
			WHEN "01110001" => U_I <= "00000001001100010011111000000";
			WHEN "01110010" => U_I <= "00000001001001000011111000000";
			WHEN "01110011" => U_I <= "00000010000001000011111000000";
			WHEN "01110100" => U_I <= "00000000000001111011111000000";
			WHEN "01110101" => U_I <= "00000001000010000011111000000";
			WHEN "01110110" => U_I <= "00000001000000000000000000000";
			when "01110111" => U_I <= "00000000000000000000000000000";
			
			
			-- 01111  RET
			WHEN "01111000" => U_I <= "00000001110111000001111000000";
			WHEN "01111001" => U_I <= "00000001111010000001111000000";
			WHEN "01111010" => U_I <= "00000001010110000001111000000";
			WHEN "01111011" => U_I <= "00000010000010000011111000000";
			WHEN "01111100" => U_I <= "00000001001000110011111000000";
			WHEN "01111101" => U_I <= "00000001111101000000000000000";
			WHEN "01111110" => U_I <= "00000000000000000000000000000";
			WHEN "01111111" => U_I <= "00000000000000000000000000000";
			
		
	      	-- 10000  MOV A,[DPTR]
			WHEN "10000000" => U_I <= "00000010000010000000010000000"; -- MAR = DPTR, RD MREQ
			WHEN "10000001" => U_I <= "00000100111000110000000000000"; -- MDR=DEX,RD MREQ,ACC=MDR,RST UPC 
			WHEN "10000010" => U_I <= "00000100011111001000000000000"; -- PC = ACC, Reset UPC
			WHEN "10000011" => U_I <= "00000000000000000000000000000";
	
			-- 10001  PUSH ACC
			WHEN "10001000" => U_I <= "00000010000100000010110000000"; -- MAR = SP
			WHEN "10001001" => U_I <= "00000001111000100001001000000"; -- MDR = ACC, WR MREQ
			WHEN "10001010" => U_I <= "00110001001001000110000000000"; -- SP++, RST UPC
			WHEN "10001011" => U_I <= "00000000000000000000000000000"; -- 
			WHEN "10001100" => U_I <= "00000000000000000000000000000"; -- 
			WHEN "10001101" => U_I <= "00000000000000000000000000000"; -- 
			WHEN "10001110" => U_I <= "00000000000000000000000000000";
			WHEN "10001111" => U_I <= "00000000000000000000000000000";

			-- 10010  POP ACC
			WHEN "10010000" => U_I <= "00000010111010000010011000000"; -- ACC = SP
			WHEN "10010001" => U_I <= "10100001001110000010011000000"; -- SP= ACC+(-1)
			WHEN "10010010" => U_I <= "00000010000100000010110000000"; -- MAR = SP
			WHEN "10010011" => U_I <= "00000100111000110000000000000"; -- MDR=DEX,RD MREQ,ACC=MDR, RST UPC
			WHEN "10010100" => U_I <= "00000000000000000000000000000"; -- 
			WHEN "10010101" => U_I <= "00000000000000000000000000000"; -- 
			WHEN "10010110" => U_I <= "00000000000000000000000000000";
			WHEN "10010111" => U_I <= "00000000000000000000000000000";

	-- 10011 ROTD A
			WHEN "10011000" => U_I <= "11000000000011000100000000000";-- para negativo
			WHEN "10011001" => U_I <= "00000000000000000000000000000";-- CONSERVAR LA BANDERA

	-- 10100 ROTD ACC
			WHEN "10100000" => U_I <= "11000000000111000100000000000";-- para negativo
			WHEN "10100001" => U_I <= "00000000000000000000000000000";-- CONSERVAR LA BANDERA

	-- 10101 PASAR ACC
			WHEN "10101000" => U_I <= "00000000000111000100000000000";-- para negativo Q-1
			WHEN "10101001" => U_I <= "00000000000000000000000000000";-- CONSERVAR LA BANDERA

	-- 10110 SUB ACC A
			WHEN "10110000" => U_I <= "00110001011011000101100000000";-- -A
			WHEN "10110001" => U_I <= "00101001111011000100000000000";-- ACC=ACC+A 
			WHEN "10110010" => U_I <= "00000000000000000000000000000";-- CONSERVAR LA BANDERA
	
		
	-- 11000 DESPL ACC
			WHEN "11000000" => U_I <= "10000001111111000100011000000";
			WHEN "11000001" => U_I <= "00000000000000000000000000000";-- DESPL ACC 
		
	-- 11001 DEC ACC
			WHEN "11001000" => U_I <= "00101001111110000100000000000";
			WHEN "11001001" => U_I <= "00000000000000000000000000000";-- DESPL ACC 
	
	-- 11010 MOV [DPTR],CTE,--- Es la unión de MOV ACC, CTE y MOV[DPTR],ACC
			WHEN "11010000" => U_I <= "00000010000000000000010000000"; -- MAR = PC, RD MREQ
			WHEN "11010001" => U_I <= "00110001000000000001000000000"; -- PC = PC + 1, RD MREQ
			WHEN "11010010" => U_I <= "00000001111000110010011000000"; -- ACC = DATA, RD MREQ, Reset UPC
			WHEN "11010011" => U_I <= "00000010000010000000010000000"; -- MAR=DPTR
			WHEN "11010100" => U_I <= "00000100000111111110000000000"; -- MDR = ACC, WR MREQ, RST UPC
			WHEN "11010101" => U_I <= "00000000000000000000000000000";	 
   --	11011 MOV DPTR,CTE
	
			WHEN "11011000" => U_I <= "00000010000000000000010000000"; -- MAR = PC, RD MREQ
			WHEN "11011001" => U_I <= "00110001000000000001000000000"; -- PC = PC + 1, RD MREQ
			WHEN "11011010" => U_I <= "00000001111000110010011000000"; -- ACC = DATA, RD MREQ, Reset UPC
			WHEN "11011011" => U_I <= "00000100000111111110000000000"; -- DPTR = ACC , Reset UPC
			WHEN "11011100" => U_I <= "00000000000000000000000000000";
	-- 11100 DEC [DPTR]
	
			WHEN "11100000" => U_I <= "00000010000010000000010000000"; -- MAR = DPTR, RD MREQ
			WHEN "11100001" => U_I <= "00000100111000110000000000000"; -- MDR=DEX,RD MREQ,ACC=MDR,RST UPC 
			WHEN "11100010" => U_I <= "00101001111110000100000000000"; -- DEC ACC
			WHEN "11100011" => U_I <= "00000010000010000000010000000"; -- MAR=DPTR
			WHEN "11100100" => U_I <= "00000100000111111110000000000"; -- MDR = ACC, WR MREQ, RST UPC
			WHEN "11100101" => U_I <= "00000000000000000000000000000";
	-- 11101 AND A,CTE
	
			WHEN "11101000" => U_I <= "00000010000000000000010000000"; -- MAR = PC, RD MREQ
			WHEN "11101001" => U_I <= "00110001000000000001000000000"; -- PC = PC + 1, RD MREQ
			WHEN "11101010" => U_I <= "00000001111000110010011000000"; -- ACC = DATA, RD MREQ, Reset UPC
			WHEN "11101011" => U_I <= "00010001111011000100011000000"; -- ACC = ACC and A, Reset UPC
			WHEN "11101100" => U_I <= "00000001111111000100000000000"; -- PC = ACC, Reset UPC
			WHEN "11101101" => U_I <= "00000000000000000000000000000";	
	
	-- 11110 MOV [DPTR],A
			
			WHEN "11110000" => U_I <= "00000001111011000101001000000"; -- ACC = A , Reset UPC
			WHEN "11110001" => U_I <= "00000010000010000000010000000"; -- MAR=DPTR
			WHEN "11110010" => U_I <= "00000100000111111110000000000"; -- MDR = ACC, WR MREQ, RST UPC
			WHEN "11110011" => U_I <= "00000000000000000000000000000";	  
   
	-- 11111 STRMEM DIR, CTE
			
			WHEN "11111000" => U_I <= "00000010000000000000010000000"; -- MAR = PC, RD MREQ
			WHEN "11111001" => U_I <= "00110001000000000001000000000"; -- PC = PC + 1, RD MREQ
			WHEN "11111010" => U_I <= "00000100000111111110000000000"; -- DPTR = DATA, RD MREQ, Reset UPC
			WHEN "11111011" => U_I <= "00000010000000000000010000000"; -- MAR = PC, RD MREQ
			WHEN "11111100" => U_I <= "00110001000000000001000000000"; -- PC = PC + 1, RD MREQ
			WHEN "11111101" => U_I <= "00000001111000110010011000000"; -- ACC = DATA, RD MREQ, Reset UPC
			WHEN "11111110" => U_I <= "00000010000010000000010000000"; -- MAR=DPTR
			WHEN "11111111" => U_I <= "00000100000111111110000000000"; -- MDR = ACC, WR MREQ, RST UPC
			

			WHEN others => U_I <= (others => 'X');
		END CASE;
	END PROCESS;
END ARCHITECTURE Behavioral;




